<ColorDecisionList>
    <ColorDecision>
        <ColorCorrection id="green">
            <SOPNode>
                <Slope>0.7 1.5 0.7</Slope>
                <Offset>-0.05 0.1 -0.05</Offset>
                <Power>1.0 0.9 1.0</Power>
            </SOPNode>
            <SatNode>
                <Saturation>1.0</Saturation>
            </SatNode>
        </ColorCorrection>
    </ColorDecision>
</ColorDecisionList>