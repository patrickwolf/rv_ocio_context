<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="HSO_0510_comp_BOT_v003">
			<SOPNode>
				<Slope>0.9163 0.9416 0.9332</Slope>
				<Offset>0.0046 -0.0018 0.0046</Offset>
				<Power>1.0131 0.9955 1.0066</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1.0000</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
