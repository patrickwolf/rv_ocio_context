<ColorDecisionList>
    <ColorDecision>
        <ColorCorrection id="red">
            <SOPNode>
                <Slope>1.5 0.7 0.7</Slope>
                <Offset>0.1 -0.05 -0.05</Offset>
                <Power>0.9 1.0 1.0</Power>
            </SOPNode>
            <SatNode>
                <Saturation>1.0</Saturation>
            </SatNode>
        </ColorCorrection>
    </ColorDecision>
</ColorDecisionList>